`timescale 10ns/1ps
module TB_ADDER;
 	reg	[31:0] A;
	reg	[31:0] B;
	wire	      C_OUT;
	wire    [31:0] SUM;

ADDER #(32) ADDER (
	.A (A),
	.B (B),
	.C_IN (1'b0),
	.SUM (SUM),
	.C_OUT (C_OUT)
);
initial begin
	A = 32'b0000_0000_0000_0000_0000_0000_1111_0001; // 241
	B = 32'b0000_0000_0000_0000_0000_0000_1011_0001; // 177
#2
	A = 32'b1100_0000_1111_0000_1111_0000_0000_0010; // -1057951742
	B = 32'b0000_0000_0000_0000_0000_0000_1111_0001;
#2
	A = 32'b1111_0000_1111_0000_1111_0000_0000_0010; // to show carryout
	B = 32'b0100_0000_0000_0000_0000_0000_1111_0001;
#2

$finish();
end

endmodule
