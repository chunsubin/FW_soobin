`timescale 10ns/1ps
module tb_dec;

wire [3:0] Dout;
reg  [1:0] Din;
reg  Enable;


 // Form : module DEC2_to_4 ([3:0] Dout,[1:0] Din,Enable);
 DEC2_to_4 mydec (
	.Dout (Dout),
	.Din  (Din),
	.Enable (Enable)
 );

 initial 
 begin
    Enable = 0; Din = 2'b01;
 #1 Enable = 0; Din = 2'b00;
 #1 Enable = 1; Din = 2'b01;
 #1 Enable = 0; Din = 2'b01;
 #1 Enable = 1; Din = 2'b11;
 #5;  // why comment
 end

endmodule

